package spi_agent_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "./../utils/config_macro.svh"
	
	`include "spi_seq_item.svh"
	`include "spi_agent_config.svh"
	`include "spi_driver.svh"
	`include "spi_monitor.svh"
	`include "spi_sequencer.svh"
	`include "spi_agent.svh"
	`include "spi_w_seq.svh"
	`include "spi_wr_seq.svh"
	`include "spi_r_seq.svh"


endpackage: spi_agent_pkg
