package spi_test_lib_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	import spi_env_pkg::*;
	import spi_agent_pkg::*;

	`include "spi_test_base.svh"
	`include "spi_wr_test.svh"
	`include "spi_w_test.svh"
	`include "spi_r_test.svh"

endpackage: spi_test_lib_pkg
