package spi_env_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	import spi_agent_pkg::*;

	`include "spi_env_config.svh"
	`include "spi_scoreboard.svh"
	`include "spi_environment.svh"

endpackage: spi_env_pkg
